module cipher

import encoding.binary

// aead_chacha20_poly1305_encrypt encrypts and authenticates data
// RFC 8439 Section 2.8
pub fn aead_chacha20_poly1305_encrypt(key []u8, nonce []u8, aad []u8, plaintext []u8) ![]u8 {
	if key.len != 32 {
		return error('invalid key length: ${key.len}, expected 32')
	}
	if nonce.len != 12 {
		return error('invalid nonce length: ${nonce.len}, expected 12')
	}
	
	// 1. Init ChaCha20 with Key and Nonce
	mut chacha := new_chacha20(key, nonce)!
	
	// 2. Generate Poly1305 Key
	// "OTK" (One-Time Key) - generated by encrypting 32 bytes of zeros with block counter 0
	mut poly_key := []u8{len: 32}
	chacha.set_counter(0)
	chacha.xor_key_stream(mut poly_key, [u8(0)].repeat(32))
	
	// 3. Encrypt Plaintext
	// ChaCha20 for encryption starts with block counter 1
	chacha.set_counter(1)
	mut ciphertext := []u8{len: plaintext.len}
	chacha.xor_key_stream(mut ciphertext, plaintext)
	
	// 4. Compute Poly1305 Tag
	// Input: AAD || pad(AAD) || Ciphertext || pad(Ciphertext) || len(AAD) || len(Ciphertext)
	mut mac := new_poly1305(poly_key)!
	
	// AAD
	mac.update(aad)
	if aad.len % 16 != 0 {
		mac.update([u8(0)].repeat(16 - (aad.len % 16)))
	}
	
	// Ciphertext
	mac.update(ciphertext)
	if ciphertext.len % 16 != 0 {
		mac.update([u8(0)].repeat(16 - (ciphertext.len % 16)))
	}
	
	// Lengths (64-bit le)
	mut len_buf := []u8{len: 16}
	binary.little_endian_put_u64(mut len_buf, u64(aad.len))
	binary.little_endian_put_u64(mut len_buf[8..], u64(ciphertext.len)) // Length of ciphertext = plaintext
	mac.update(len_buf)
	
	tag := mac.finish()
	
	// Result: Ciphertext || Tag
	mut result := ciphertext.clone()
	result << tag
	return result
}

// aead_chacha20_poly1305_decrypt decrypts and verifies data
pub fn aead_chacha20_poly1305_decrypt(key []u8, nonce []u8, aad []u8, ciphertext_and_tag []u8) ![]u8 {
	if key.len != 32 {
		return error('invalid key length')
	}
	if nonce.len != 12 {
		return error('invalid nonce length')
	}
	if ciphertext_and_tag.len < 16 {
		return error('ciphertext too short')
	}
	
	ciphertext := ciphertext_and_tag[..ciphertext_and_tag.len - 16]
	tag := ciphertext_and_tag[ciphertext_and_tag.len - 16..]
	
	// 1. Init ChaCha20
	mut chacha := new_chacha20(key, nonce)!
	
	// 2. Generate Poly1305 Key
	mut poly_key := []u8{len: 32}
	chacha.set_counter(0)
	chacha.xor_key_stream(mut poly_key, [u8(0)].repeat(32))
	
	// 3. Verify Tag
	mut mac := new_poly1305(poly_key)!
	
	mac.update(aad)
	if aad.len % 16 != 0 {
		mac.update([u8(0)].repeat(16 - (aad.len % 16)))
	}
	
	mac.update(ciphertext)
	if ciphertext.len % 16 != 0 {
		mac.update([u8(0)].repeat(16 - (ciphertext.len % 16)))
	}
	
	mut len_buf := []u8{len: 16}
	binary.little_endian_put_u64(mut len_buf, u64(aad.len))
	binary.little_endian_put_u64(mut len_buf[8..], u64(ciphertext.len))
	mac.update(len_buf)
	
	calc_tag := mac.finish()
	
	if !constant_time_compare(calc_tag, tag) {
		return error('poly1305 tag verification failed')
	}
	
	// 4. Decrypt
	chacha.set_counter(1)
	mut plaintext := []u8{len: ciphertext.len}
	chacha.xor_key_stream(mut plaintext, ciphertext)
	
	return plaintext
}

fn constant_time_compare(a []u8, b []u8) bool {
	if a.len != b.len { return false }
	mut res := u8(0)
	for i in 0 .. a.len {
		res |= a[i] ^ b[i]
	}
	return res == 0
}
