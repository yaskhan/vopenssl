module ecc

fn test_x25519_basepoint() {
	// Basepoint multiplication test
	// scalar = 1
	mut scalar := []u8{len: 32, init: 0}
	scalar[0] = 1
	
	mut basepoint := []u8{len: 32, init: 0}
	basepoint[0] = 9
	
	res := x25519_scalarmult_impl(scalar, basepoint)
	
	// If scalar is 1, result should be basepoint 9
	assert res[0] == 9
	for i in 1 .. 32 {
		assert res[i] == 0
	}
}

fn test_x25519_rfc7748_test_vector_1() {
	// Alice's private key, a:
	// 77076d0a7318a57d3c16c17251b26645df4c2f87ebc0992ab177fba51db92c1c
	alice_priv := [u8(0x77), 0x07, 0x6d, 0x0a, 0x73, 0x18, 0xa5, 0x7d, 0x3c, 0x16, 0xc1, 0x72, 0x51, 0xb2, 0x66, 0x45, 0xdf, 0x4c, 0x2f, 0x87, 0xeb, 0xc0, 0x99, 0x2a, 0xb1, 0x77, 0xfb, 0xa5, 0x1d, 0xb9, 0x2c, 0x1c]
	
	// Alice's public key, X25519(a, 9):
	// 8520f0098930a754748b7ddcb43ef75a0dbf3a0d26381af4eba4a98eaa9b4e6a
	
	basepoint := []u8{len: 32, init: 0}
	basepoint[0] = 9
	
	res := x25519_scalarmult_impl(alice_priv, basepoint)
	
	expected := [u8(0x85), 0x20, 0xf0, 0x09, 0x89, 0x30, 0xa7, 0x54, 0x74, 0x8b, 0x7d, 0xdc, 0xb4, 0x3e, 0xf7, 0x5a, 0x0d, 0xbf, 0x3a, 0x0d, 0x26, 0x38, 0x1a, 0xf4, 0xeb, 0xa4, 0xa9, 0x8e, 0xaa, 0x9b, 0x4e, 0x6a]
	
	for i in 0 .. 32 {
		assert res[i] == expected[i]
	}
}
