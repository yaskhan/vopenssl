module tls

// TLS protocol versions
pub const version_tls_10 = u16(0x0301)
pub const version_tls_11 = u16(0x0302)
pub const version_tls_12 = u16(0x0303)
pub const version_tls_13 = u16(0x0304)

// TLS content types (record layer)
pub const content_type_change_cipher_spec = u8(20)
pub const content_type_alert = u8(21)
pub const content_type_handshake = u8(22)
pub const content_type_application_data = u8(23)

// TLS handshake message types
pub const handshake_type_hello_request = u8(0)
pub const handshake_type_client_hello = u8(1)
pub const handshake_type_server_hello = u8(2)
pub const handshake_type_new_session_ticket = u8(4)
pub const handshake_type_end_of_early_data = u8(5)
pub const handshake_type_encrypted_extensions = u8(8)
pub const handshake_type_certificate = u8(11)
pub const handshake_type_server_key_exchange = u8(12)
pub const handshake_type_certificate_request = u8(13)
pub const handshake_type_server_hello_done = u8(14)
pub const handshake_type_certificate_verify = u8(15)
pub const handshake_type_client_key_exchange = u8(16)
pub const handshake_type_finished = u8(20)
pub const handshake_type_key_update = u8(24)
pub const handshake_type_message_hash = u8(254)

// TLS alert levels
pub const alert_level_warning = u8(1)
pub const alert_level_fatal = u8(2)

// TLS alert descriptions
pub const alert_close_notify = u8(0)
pub const alert_unexpected_message = u8(10)
pub const alert_bad_record_mac = u8(20)
pub const alert_decryption_failed = u8(21)
pub const alert_record_overflow = u8(22)
pub const alert_decompression_failure = u8(30)
pub const alert_handshake_failure = u8(40)
pub const alert_no_certificate = u8(41)
pub const alert_bad_certificate = u8(42)
pub const alert_unsupported_certificate = u8(43)
pub const alert_certificate_revoked = u8(44)
pub const alert_certificate_expired = u8(45)
pub const alert_certificate_unknown = u8(46)
pub const alert_illegal_parameter = u8(47)
pub const alert_unknown_ca = u8(48)
pub const alert_access_denied = u8(49)
pub const alert_decode_error = u8(50)
pub const alert_decrypt_error = u8(51)
pub const alert_export_restriction = u8(60)
pub const alert_protocol_version = u8(70)
pub const alert_insufficient_security = u8(71)
pub const alert_internal_error = u8(80)
pub const alert_inappropriate_fallback = u8(86)
pub const alert_user_canceled = u8(90)
pub const alert_no_renegotiation = u8(100)
pub const alert_missing_extension = u8(109)
pub const alert_unsupported_extension = u8(110)
pub const alert_certificate_unobtainable = u8(111)
pub const alert_unrecognized_name = u8(112)
pub const alert_bad_certificate_status_response = u8(113)
pub const alert_bad_certificate_hash_value = u8(114)
pub const alert_unknown_psk_identity = u8(115)
pub const alert_certificate_required = u8(116)
pub const alert_no_application_protocol = u8(120)

// TLS extension types
pub const extension_server_name = u16(0)
pub const extension_max_fragment_length = u16(1)
pub const extension_status_request = u16(5)
pub const extension_supported_groups = u16(10)
pub const extension_ec_point_formats = u16(11)
pub const extension_signature_algorithms = u16(13)
pub const extension_use_srtp = u16(14)
pub const extension_heartbeat = u16(15)
pub const extension_alpn = u16(16)
pub const extension_signed_certificate_timestamp = u16(18)
pub const extension_client_certificate_type = u16(19)
pub const extension_server_certificate_type = u16(20)
pub const extension_padding = u16(21)
pub const extension_encrypt_then_mac = u16(22)
pub const extension_extended_master_secret = u16(23)
pub const extension_session_ticket = u16(35)
pub const extension_pre_shared_key = u16(41)
pub const extension_early_data = u16(42)
pub const extension_supported_versions = u16(43)
pub const extension_cookie = u16(44)
pub const extension_psk_key_exchange_modes = u16(45)
pub const extension_certificate_authorities = u16(47)
pub const extension_oid_filters = u16(48)
pub const extension_post_handshake_auth = u16(49)
pub const extension_signature_algorithms_cert = u16(50)
pub const extension_key_share = u16(51)
pub const extension_renegotiation_info = u16(0xff01)

// Supported groups (curves)
pub const supported_group_secp256r1 = u16(23)
pub const supported_group_secp384r1 = u16(24)
pub const supported_group_secp521r1 = u16(25)
pub const supported_group_x25519 = u16(29)
pub const supported_group_x448 = u16(30)

// EC point formats
pub const ec_point_format_uncompressed = u8(0)
pub const ec_point_format_ansix962_compressed_prime = u8(1)
pub const ec_point_format_ansix962_compressed_char2 = u8(2)

// Signature algorithms
pub const signature_rsa_pkcs1_sha256 = u16(0x0401)
pub const signature_rsa_pkcs1_sha384 = u16(0x0501)
pub const signature_rsa_pkcs1_sha512 = u16(0x0601)
pub const signature_ecdsa_secp256r1_sha256 = u16(0x0403)
pub const signature_ecdsa_secp384r1_sha384 = u16(0x0503)
pub const signature_ecdsa_secp521r1_sha512 = u16(0x0603)
pub const signature_rsa_pss_rsae_sha256 = u16(0x0804)
pub const signature_rsa_pss_rsae_sha384 = u16(0x0805)
pub const signature_rsa_pss_rsae_sha512 = u16(0x0806)
pub const signature_ed25519 = u16(0x0807)
pub const signature_ed448 = u16(0x0808)
pub const signature_rsa_pss_pss_sha256 = u16(0x0809)
pub const signature_rsa_pss_pss_sha384 = u16(0x080a)
pub const signature_rsa_pss_pss_sha512 = u16(0x080b)
pub const signature_rsa_pkcs1_sha1 = u16(0x0201)
pub const signature_ecdsa_sha1 = u16(0x0203)

// TLS record size limits
pub const max_plaintext_length = 16384 // 2^14 bytes

pub const max_ciphertext_length = 16384 + 2048 // plaintext + expansion

pub const max_handshake_length = 65536 // maximum handshake message size
