module main

fn main() {
	mut h0 := u32(0x6a09e667)
	mut h1 := u32(0xbb67ae85)
	mut h2 := u32(0x3c6ef372)
	mut h3 := u32(0xa54ff53a)
	mut h4 := u32(0x510e527f)
	mut h5 := u32(0x9b05688c)
	mut h6 := u32(0x1f83d9ab)
	mut h7 := u32(0x5be0cd19)

	k := [
		u32(0x428a2f98), 0x71374491, 0xb5c0fbcf, 0xe9b5dba5, 0x3956c25b, 0x59f111f1, 0x923f82a4, 0xab1c5ed5,
		0xd807aa98, 0x12835b01, 0x243185be, 0x550c7dc3, 0x72be5d74, 0x80deb1fe, 0x9bdc06a7, 0xc19bf174,
		0xe49b69c1, 0xefbe4786, 0x0fc19dc6, 0x240ca1cc, 0x2de92c6f, 0x4a7484aa, 0x5cb0a9dc, 0x76f988da,
		0x983e5152, 0xa831c66d, 0xb00327c8, 0xbf597fc7, 0xc6e00bf3, 0xd5a79147, 0x06ca6351, 0x14292967,
		0x27b70a85, 0x2e1b2138, 0x4d2c6dfc, 0x53380d13, 0x650a7354, 0x766a0abb, 0x81c2c92e, 0x92722c85,
		0xa2bfe8a1, 0xa81a664b, 0xc24b8b70, 0xc76c51a3, 0xd192e819, 0xd6990624, 0xf40e3585, 0x106aa070,
		0x19a4c116, 0x1e376c08, 0x2748774c, 0x34b0bcb5, 0x391c0cb3, 0x4ed8aa4a, 0x5b9cca4f, 0x682e6ff3,
		0x748f82ee, 0x78a5636f, 0x84c87814, 0x8cc70208, 0x90befffa, 0xa4506ceb, 0xbef9a3f7, 0xc67178f2,
	]

	// Block for empty string: 80 00 ... 00
	mut w := [64]u32{}
	w[0] = 0x80000000
	// 1..15 are 0
	
	// Extend
	for i in 16 .. 64 {
		s0 := (w[i-15] >> 7 | w[i-15] << 25) ^ (w[i-15] >> 18 | w[i-15] << 14) ^ (w[i-15] >> 3)
		s1 := (w[i-2] >> 17 | w[i-2] << 15) ^ (w[i-2] >> 19 | w[i-2] << 13) ^ (w[i-2] >> 10)
		w[i] = w[i-16] + s0 + w[i-7] + s1
	}
	
	mut a := h0
	mut b := h1
	mut c := h2
	mut d := h3
	mut e := h4
	mut f := h5
	mut g := h6
	mut h := h7
	
	for i in 0 .. 64 {
		s1 := (e >> 6 | e << 26) ^ (e >> 11 | e << 21) ^ (e >> 25 | e << 7)
		ch := (e & f) ^ ((~e) & g)
		temp1 := h + s1 + ch + k[i] + w[i]
		s0 := (a >> 2 | a << 30) ^ (a >> 13 | a << 19) ^ (a >> 22 | a << 10)
		maj := (a & b) ^ (a & c) ^ (b & c)
		temp2 := s0 + maj
		
		h = g
		g = f
		f = e
		e = d + temp1
		d = c
		c = b
		b = a
		a = temp1 + temp2
	}
	
	h0 += a
	h1 += b
	h2 += c
	h3 += d
	h4 += e
	h5 += f
	h6 += g
	h7 += h
	
	println('${h0:08x}${h1:08x}${h2:08x}${h3:08x}${h4:08x}${h5:08x}${h6:08x}${h7:08x}')
}
